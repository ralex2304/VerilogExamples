bind fifo fifo_assertions fifo_assertions_inst (.*);
